VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_timer
  CLASS BLOCK ;
  FOREIGN user_proj_timer ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 3000.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2934.920 4.000 2935.520 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END io_in[10]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2665.640 4.000 2666.240 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2396.360 4.000 2396.960 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2127.080 4.000 2127.680 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1857.800 4.000 1858.400 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1588.520 4.000 1589.120 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1319.240 4.000 1319.840 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1049.960 4.000 1050.560 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 780.680 4.000 781.280 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 511.400 4.000 512.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2755.400 4.000 2756.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END io_oeb[10]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2486.120 4.000 2486.720 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2216.840 4.000 2217.440 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1947.560 4.000 1948.160 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1678.280 4.000 1678.880 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1409.000 4.000 1409.600 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1139.720 4.000 1140.320 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 870.440 4.000 871.040 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.160 4.000 601.760 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2845.160 4.000 2845.760 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END io_out[10]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2575.880 4.000 2576.480 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2306.600 4.000 2307.200 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2037.320 4.000 2037.920 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1768.040 4.000 1768.640 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1498.760 4.000 1499.360 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1229.480 4.000 1230.080 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 960.200 4.000 960.800 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.920 4.000 691.520 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END io_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 2986.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 2986.800 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END wb_rst_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 2986.645 ;
      LAYER met1 ;
        RECT 4.670 10.640 194.120 2986.800 ;
      LAYER met2 ;
        RECT 4.690 4.280 176.210 2986.745 ;
        RECT 4.690 4.000 49.490 4.280 ;
        RECT 50.330 4.000 149.310 4.280 ;
        RECT 150.150 4.000 176.210 4.280 ;
      LAYER met3 ;
        RECT 4.000 2935.920 176.230 2986.725 ;
        RECT 4.400 2934.520 176.230 2935.920 ;
        RECT 4.000 2846.160 176.230 2934.520 ;
        RECT 4.400 2844.760 176.230 2846.160 ;
        RECT 4.000 2756.400 176.230 2844.760 ;
        RECT 4.400 2755.000 176.230 2756.400 ;
        RECT 4.000 2666.640 176.230 2755.000 ;
        RECT 4.400 2665.240 176.230 2666.640 ;
        RECT 4.000 2576.880 176.230 2665.240 ;
        RECT 4.400 2575.480 176.230 2576.880 ;
        RECT 4.000 2487.120 176.230 2575.480 ;
        RECT 4.400 2485.720 176.230 2487.120 ;
        RECT 4.000 2397.360 176.230 2485.720 ;
        RECT 4.400 2395.960 176.230 2397.360 ;
        RECT 4.000 2307.600 176.230 2395.960 ;
        RECT 4.400 2306.200 176.230 2307.600 ;
        RECT 4.000 2217.840 176.230 2306.200 ;
        RECT 4.400 2216.440 176.230 2217.840 ;
        RECT 4.000 2128.080 176.230 2216.440 ;
        RECT 4.400 2126.680 176.230 2128.080 ;
        RECT 4.000 2038.320 176.230 2126.680 ;
        RECT 4.400 2036.920 176.230 2038.320 ;
        RECT 4.000 1948.560 176.230 2036.920 ;
        RECT 4.400 1947.160 176.230 1948.560 ;
        RECT 4.000 1858.800 176.230 1947.160 ;
        RECT 4.400 1857.400 176.230 1858.800 ;
        RECT 4.000 1769.040 176.230 1857.400 ;
        RECT 4.400 1767.640 176.230 1769.040 ;
        RECT 4.000 1679.280 176.230 1767.640 ;
        RECT 4.400 1677.880 176.230 1679.280 ;
        RECT 4.000 1589.520 176.230 1677.880 ;
        RECT 4.400 1588.120 176.230 1589.520 ;
        RECT 4.000 1499.760 176.230 1588.120 ;
        RECT 4.400 1498.360 176.230 1499.760 ;
        RECT 4.000 1410.000 176.230 1498.360 ;
        RECT 4.400 1408.600 176.230 1410.000 ;
        RECT 4.000 1320.240 176.230 1408.600 ;
        RECT 4.400 1318.840 176.230 1320.240 ;
        RECT 4.000 1230.480 176.230 1318.840 ;
        RECT 4.400 1229.080 176.230 1230.480 ;
        RECT 4.000 1140.720 176.230 1229.080 ;
        RECT 4.400 1139.320 176.230 1140.720 ;
        RECT 4.000 1050.960 176.230 1139.320 ;
        RECT 4.400 1049.560 176.230 1050.960 ;
        RECT 4.000 961.200 176.230 1049.560 ;
        RECT 4.400 959.800 176.230 961.200 ;
        RECT 4.000 871.440 176.230 959.800 ;
        RECT 4.400 870.040 176.230 871.440 ;
        RECT 4.000 781.680 176.230 870.040 ;
        RECT 4.400 780.280 176.230 781.680 ;
        RECT 4.000 691.920 176.230 780.280 ;
        RECT 4.400 690.520 176.230 691.920 ;
        RECT 4.000 602.160 176.230 690.520 ;
        RECT 4.400 600.760 176.230 602.160 ;
        RECT 4.000 512.400 176.230 600.760 ;
        RECT 4.400 511.000 176.230 512.400 ;
        RECT 4.000 422.640 176.230 511.000 ;
        RECT 4.400 421.240 176.230 422.640 ;
        RECT 4.000 332.880 176.230 421.240 ;
        RECT 4.400 331.480 176.230 332.880 ;
        RECT 4.000 243.120 176.230 331.480 ;
        RECT 4.400 241.720 176.230 243.120 ;
        RECT 4.000 153.360 176.230 241.720 ;
        RECT 4.400 151.960 176.230 153.360 ;
        RECT 4.000 63.600 176.230 151.960 ;
        RECT 4.400 62.200 176.230 63.600 ;
        RECT 4.000 10.715 176.230 62.200 ;
      LAYER met4 ;
        RECT 24.215 17.175 47.545 916.465 ;
  END
END user_proj_timer
END LIBRARY

